

////////////////////////////////////////////////////////////////////////////////
// 
// N-BIT DEMUX
//
////////////////////////////////////////////////////////////////////////////////
module demux (
    bits_out, sel, bit_in
);
    parameter SEL_BITS = 1;
    output [2**SEL_BITS - 1: 0] bits_out;
    input [SEL_BITS-1:0] sel;
    input bit_in;
    
    assign bits_out = (bit_in << sel);
endmodule

////////////////////////////////////////////////////////////////////////////////
// 
// N-BIT MUX
//
////////////////////////////////////////////////////////////////////////////////
module mux (
    out, sel, bits_in
);
    parameter SEL_BITS = 1;
    output out;
    input [SEL_BITS-1:0] sel;
    input [2**SEL_BITS - 1: 0] bits_in;

    assign out = bits_in[sel];
endmodule
