///////////////////////////////////////////////////////////////////////////////
// 
// N-BIT ADDER
//
///////////////////////////////////////////////////////////////////////////////
module adder(sum, cout, a, b, cin);

parameter BITS = 16;

output [BITS-1:0] sum;
output cout;

input [BITS-1:0] a;
input [BITS-1:0] b;
input cin;

assign {cout, sum} = a + b + cin;

endmodule